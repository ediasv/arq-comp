library ieee;
use ieee.std_logic_1164.all;
ieee.numeric_std.all
