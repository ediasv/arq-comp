library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity rom is
  port (clk      : in  std_logic;
        endereco : in  unsigned(6 downto 0);
        dado     : out unsigned(14 downto 0)
       );
end entity;

--TAMANHO DA INSTRUÇÃO: 15 bits
--ROM síncrona de 128 enderecos

architecture a_rom of rom is
  type mem is array (0 to 127) of unsigned(14 downto 0);
  constant conteudo_rom : mem := (
    0      => "000100000100101", -- LD R1, 2
    1      => "001001000000101", -- LD R2, 32
    2      => "011100000010101", -- LD R7, 1
    3      => "000100000010100", -- MV ACC, R1
    4      => "000100000011011", -- SW ACC, R1
    5      => "000100001110001", -- ADD ACC, R7
    6      => "000000110000100", -- MV R1, ACC
    7      => "000100000100100", -- MV ACC, R2
    8      => "000100000010010", -- SUB ACC, R1
    9      => "000000000100111", -- BEQ 2
    10     => "000000000110110", -- JMP 3
    11     => "000000000000000", -- NOP
    others => (others => '0')
  );

  signal dado_sig : unsigned(14 downto 0) := conteudo_rom(0);
begin
  process (clk)
  begin
    if (rising_edge(clk)) then
      if (endereco >= 0 and endereco <= 127) then
        dado_sig <= conteudo_rom(to_integer(endereco));
      else
        dado_sig <= (others => '0');
      end if;
    end if;
  end process;

  dado <= dado_sig;
end architecture;
